module add(
  inout a,
  input b,
  output c
);
  assign c = a^b;
endmodule
